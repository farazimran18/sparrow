package yarp_pkg;

endpackage
