import yarp_pkg::*;

module yarp_branch_control (
    // Source operands
    input logic [31:0] opr_a_i,
    input logic [31:0] opr_b_i,

    // Branch Type
    input logic       is_b_type_ctl_i,
    input logic [2:0] instr_func3_ctl_i,

    // Branch outcome
    output logic branch_taken_o
  );

  // Write your logic here...

endmodule
