package yarp_pkg;

  localparam int XLEN = 32;

endpackage
